module main

struct Post {
	date string
	estimated_read_time_minutes int
	content string
}
